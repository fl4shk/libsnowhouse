../../../../hw/verilog/LcvMulAcc.sv