../../submodules/libcheesevoyage/hw/verilog/LcvMulAcc.sv